CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 250 30 120 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
72
8 SPDT PB~
217 300 689 0 10 18
0 4 4 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
5 RESET
-14 -15 21 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
5305 0 0
2
44316.3 0
0
10 3-In NAND~
219 428 863 0 4 22
0 8 4 9 28
0
0 0 112 0
5 74F10
-18 -28 17 -20
4 U28A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 21 0
1 U
34 0 0
2
5.89983e-315 0
0
9 2-In NOR~
219 2117 1306 0 3 22
0 7 6 5
0
0 0 112 0
6 74LS02
-21 -24 21 -16
4 U29A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 22 0
1 U
969 0 0
2
44316.3 1
0
9 Inverter~
13 2070 1314 0 2 22
0 4 6
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U10E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 10 0
1 U
8402 0 0
2
44316.3 2
0
14 NO PushButton~
191 297 751 0 2 5
0 27 2
0
0 0 4720 0
0
6 ANSWER
-21 -20 21 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3751 0 0
2
5.89983e-315 0
0
5 7474~
219 1510 426 0 6 22
0 4 42 38 4 96 33
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U27B
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 20 0
1 U
4292 0 0
2
44316.3 4
0
5 7474~
219 1583 425 0 6 22
0 4 41 38 4 97 32
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U27A
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 20 0
1 U
6118 0 0
2
44316.3 5
0
5 7474~
219 1653 425 0 6 22
0 4 40 38 4 98 31
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U26B
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 19 0
1 U
34 0 0
2
44316.3 6
0
5 7474~
219 1726 425 0 6 22
0 4 39 38 4 99 30
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U26A
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 19 0
1 U
6357 0 0
2
44316.3 7
0
7 74LS157
122 1460 288 0 14 29
0 29 14 30 13 31 12 32 11 33
2 39 40 41 42
0
0 0 4336 270
6 74F157
-21 -60 21 -52
3 U25
51 0 72 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
319 0 0
2
44316.3 8
0
7 Ground~
168 1414 247 0 1 3
0 2
0
0 0 53360 180
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3976 0 0
2
44316.3 9
0
7 Ground~
168 909 247 0 1 3
0 2
0
0 0 53360 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7634 0 0
2
44316.3 10
0
7 74LS157
122 955 288 0 14 29
0 29 18 34 17 35 16 36 15 37
2 43 44 45 46
0
0 0 4336 270
6 74F157
-21 -60 21 -52
3 U24
51 0 72 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
523 0 0
2
44316.3 11
0
5 7474~
219 1221 425 0 6 22
0 4 43 38 4 100 34
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U23B
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 18 0
1 U
6748 0 0
2
44316.3 12
0
5 7474~
219 1148 425 0 6 22
0 4 44 38 4 101 35
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U23A
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 18 0
1 U
6901 0 0
2
44316.3 13
0
5 7474~
219 1078 425 0 6 22
0 4 45 102 4 103 36
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U22B
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 17 0
1 U
842 0 0
2
44316.3 14
0
5 7474~
219 1005 426 0 6 22
0 4 46 38 4 104 37
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U22A
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 17 0
1 U
3277 0 0
2
44316.3 15
0
12 Hex Display~
7 695 383 0 16 19
10 30 31 32 33 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
3 LSB
-11 -38 10 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4212 0 0
2
44316.3 16
0
12 Hex Display~
7 610 384 0 16 19
10 34 35 36 37 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
3 MSB
-11 -38 10 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4720 0 0
2
44316.3 17
0
8 Hex Key~
166 373 377 0 11 12
0 26 25 24 23 0 0 0 0 0
0 48
0
0 0 4656 0
0
2 IA
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5551 0 0
2
44316.3 18
0
5 7474~
219 1772 954 0 6 22
0 4 92 38 4 105 48
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
6986 0 0
2
44316.3 19
0
5 7474~
219 1846 960 0 6 22
0 4 91 38 4 106 49
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
8745 0 0
2
44316.3 20
0
5 7474~
219 1916 960 0 6 22
0 4 90 38 4 107 50
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
9592 0 0
2
44316.3 21
0
5 7474~
219 1989 960 0 6 22
0 4 89 38 4 108 51
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U3B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 3 0
1 U
8748 0 0
2
44316.3 22
0
7 Ground~
168 1735 781 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
44316.3 23
0
9 2-In XOR~
219 2157 1069 0 3 22
0 51 82 93
0
0 0 112 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
631 0 0
2
44316.3 24
0
10 2-In NAND~
219 2244 1128 0 3 22
0 51 82 95
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9466 0 0
2
44316.3 25
0
10 2-In NAND~
219 2311 1151 0 3 22
0 95 94 58
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3266 0 0
2
44316.3 26
0
9 2-In XOR~
219 2299 1078 0 3 22
0 93 52 81
0
0 0 112 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7693 0 0
2
44316.3 27
0
10 2-In NAND~
219 2245 1175 0 3 22
0 93 52 94
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3723 0 0
2
44316.3 28
0
5 7474~
219 2260 1263 0 6 22
0 4 59 38 5 109 52
0
0 0 4208 512
4 7474
7 -60 35 -52
3 U5A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 5 0
1 U
3440 0 0
2
44316.3 29
0
5 7474~
219 1353 962 0 6 22
0 4 67 64 4 110 69
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U5B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 5 0
1 U
6263 0 0
2
44316.3 30
0
4 4539
219 1808 828 0 14 29
0 49 48 16 49 2 48 81 15 48
2 53 7 92 91
0
0 0 4336 270
4 4539
-14 -60 14 -52
3 U17
62 9 83 17
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
4900 0 0
2
44316.3 31
0
4 4539
219 1947 828 0 14 29
0 51 50 18 51 2 50 49 17 50
2 53 7 90 89
0
0 0 4336 270
4 4539
-14 -60 14 -52
3 U13
62 9 83 17
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
8783 0 0
2
44316.3 32
0
4 4539
219 1946 1129 0 14 29
0 82 83 14 82 2 83 72 13 83
2 53 7 86 85
0
0 0 4336 270
4 4539
-14 -60 14 -52
3 U12
62 9 83 17
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
3221 0 0
2
44316.3 33
0
4 4539
219 1808 1129 0 14 29
0 72 84 12 72 2 84 2 11 84
2 53 7 88 87
0
0 0 4336 270
4 4539
-14 -60 14 -52
3 U11
62 9 83 17
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
3215 0 0
2
44316.3 34
0
7 Ground~
168 1735 1082 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7903 0 0
2
44316.3 35
0
5 7474~
219 1989 1261 0 6 22
0 4 85 38 4 111 82
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U6A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 6 0
1 U
7121 0 0
2
44316.3 36
0
5 7474~
219 1916 1261 0 6 22
0 4 86 38 4 112 83
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U6B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 6 0
1 U
4484 0 0
2
44316.3 37
0
5 7474~
219 1846 1261 0 6 22
0 4 87 38 4 113 72
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U7A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 7 0
1 U
5996 0 0
2
44316.3 38
0
5 7474~
219 1773 1262 0 6 22
0 4 88 38 4 114 84
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U7B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 7 0
1 U
7804 0 0
2
44316.3 39
0
8 Hex Key~
166 454 376 0 11 12
0 19 20 21 22 0 0 0 0 0
0 48
0
0 0 4656 0
0
2 IB
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5523 0 0
2
44316.3 40
0
5 7474~
219 1266 963 0 6 22
0 4 71 64 4 66 63
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U8A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 8 0
1 U
3330 0 0
2
44316.3 41
0
9 2-In AND~
219 714 1067 0 3 22
0 73 53 74
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3465 0 0
2
44316.3 42
0
9 Inverter~
13 649 722 0 2 22
0 54 73
0
0 0 112 180
6 74LS04
-21 -19 21 -11
4 U10A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
8396 0 0
2
44316.3 43
0
8 2-In OR~
219 787 1048 0 3 22
0 7 74 75
0
0 0 112 0
6 74LS32
-21 -24 21 -16
4 U14A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3685 0 0
2
44316.3 44
0
9 2-In AND~
219 780 1135 0 3 22
0 53 54 55
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
7849 0 0
2
44316.3 45
0
9 2-In AND~
219 1039 1061 0 3 22
0 53 56 64
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
6343 0 0
2
44316.3 46
0
7 Pulser~
4 310 1200 0 10 12
0 115 116 56 38 0 0 5 5 2
8
0
0 0 4656 0
0
3 CLK
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7376 0 0
2
44316.3 47
0
2 +V
167 279 1011 0 1 3
0 4
0
0 0 54128 0
2 5V
-8 -22 6 -14
3 VDD
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9156 0 0
2
44316.3 48
0
5 7474~
219 863 844 0 6 22
0 4 77 56 4 117 78
0
0 0 4208 0
4 7474
7 -60 35 -52
3 U8B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 8 0
1 U
5776 0 0
2
44316.3 49
0
5 7474~
219 863 962 0 6 22
0 4 80 56 4 10 7
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U15A
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 12 0
1 U
7207 0 0
2
44316.3 50
0
5 7474~
219 866 1084 0 6 22
0 4 75 56 4 9 53
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U15B
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 12 0
1 U
4459 0 0
2
44316.3 51
0
9 2-In AND~
219 771 816 0 3 22
0 79 78 76
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
3760 0 0
2
44316.3 52
0
9 2-In AND~
219 773 926 0 3 22
0 78 8 80
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
754 0 0
2
44316.3 53
0
9 Inverter~
13 706 807 0 2 22
0 8 79
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U10B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
9767 0 0
2
44316.3 54
0
8 2-In OR~
219 804 808 0 3 22
0 29 76 77
0
0 0 112 0
6 74LS32
-21 -24 21 -16
4 U14B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
7978 0 0
2
44316.3 55
0
9 2-In AND~
219 1225 722 0 3 22
0 63 62 54
0
0 0 112 180
6 74LS08
-21 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
3142 0 0
2
44316.3 56
0
5 7474~
219 1436 962 0 6 22
0 4 65 64 4 62 70
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U18A
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 14 0
1 U
3284 0 0
2
44316.3 57
0
9 3-In AND~
219 1198 927 0 4 22
0 70 69 66 71
0
0 0 112 0
5 74F11
-18 -28 17 -20
4 U19A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 15 0
1 U
659 0 0
2
44316.3 58
0
9 2-In XOR~
219 1381 1034 0 3 22
0 70 69 68
0
0 0 112 180
6 74LS86
-21 -24 21 -16
3 U1D
-2 -25 19 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3800 0 0
2
44316.3 59
0
9 2-In AND~
219 1312 1010 0 3 22
0 66 68 67
0
0 0 112 90
6 74LS08
-21 -24 21 -16
4 U16C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
6792 0 0
2
44316.3 60
0
9 2-In AND~
219 1445 1002 0 3 22
0 66 62 65
0
0 0 112 180
6 74LS08
-21 -24 21 -16
4 U16D
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
3701 0 0
2
44316.3 61
0
9 2-In AND~
219 2422 1188 0 3 22
0 53 58 61
0
0 0 112 180
6 74LS08
-21 -24 21 -16
4 U20A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
6316 0 0
2
44316.3 62
0
9 2-In AND~
219 2419 1268 0 3 22
0 52 57 60
0
0 0 112 180
6 74LS08
-21 -24 21 -16
4 U20B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
8734 0 0
2
44316.3 63
0
8 2-In OR~
219 2361 1227 0 3 22
0 60 61 59
0
0 0 112 180
6 74LS32
-21 -24 21 -16
4 U14C
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
7988 0 0
2
44316.3 64
0
9 Inverter~
13 2450 1227 0 2 22
0 53 57
0
0 0 112 270
6 74LS04
-21 -19 21 -11
4 U10C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
3217 0 0
2
44316.3 65
0
5 7474~
219 866 1171 0 6 22
0 4 55 56 4 47 29
0
0 0 4208 0
4 7474
7 -60 35 -52
4 U18B
19 -61 47 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 14 0
1 U
3965 0 0
2
44316.3 66
0
7 74LS244
143 2282 895 0 18 37
0 2 2 2 52 48 49 50 51 15
16 17 18 11 12 13 14 47 47
0
0 0 4336 0
7 74LS244
-24 -60 25 -52
3 U21
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 0 0 0
1 U
8239 0 0
2
44316.3 67
0
7 Ground~
168 273 793 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
828 0 0
2
44316.3 68
0
10 2-In NAND~
219 428 767 0 3 22
0 27 28 8
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
6187 0 0
2
44316.3 69
0
7 74LS244
143 410 473 0 18 37
0 19 20 21 22 26 25 24 23 14
13 12 11 18 17 16 15 10 10
0
0 0 4336 270
7 74LS244
-24 -60 25 -52
3 U30
53 0 74 8
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 0 0 0
1 U
7107 0 0
2
44316.3 70
0
266
2 1 4 0 0 8192 3 1 50 0 0 4
283 689
258 689
258 1020
279 1020
3 0 2 0 0 12288 0 1 0 0 41 4
283 703
283 701
273 701
273 759
2 0 4 0 0 4096 0 2 0 0 10 2
404 863
346 863
3 0 5 0 0 0 0 3 0 0 8 2
2156 1306
2156 1306
0 1 4 0 0 8192 0 0 4 225 0 3
1989 1279
1989 1314
2055 1314
2 2 6 0 0 8320 0 4 3 0 0 3
2091 1314
2091 1315
2104 1315
0 1 7 0 0 4096 0 0 3 197 0 4
1636 1029
2085 1029
2085 1297
2104 1297
0 4 5 0 0 4224 0 0 31 0 0 5
2153 1306
2265 1306
2265 1278
2266 1278
2266 1275
0 1 8 0 0 12416 0 0 56 42 0 4
501 808
559 808
559 807
691 807
1 0 4 0 0 8208 0 1 0 0 128 5
322 689
346 689
346 1254
618 1254
618 1253
0 4 4 0 0 0 0 0 68 128 0 4
865 1253
865 1254
866 1254
866 1183
5 3 9 0 0 12416 0 53 2 0 0 6
896 1066
909 1066
909 1005
388 1005
388 872
404 872
5 0 10 0 0 12416 0 52 0 0 15 6
893 944
921 944
921 620
499 620
499 436
445 436
2 0 8 0 0 0 0 55 0 0 9 3
749 935
654 935
654 807
17 18 10 0 0 0 0 72 72 0 0 4
445 440
445 436
400 436
400 440
8 3 11 0 0 12416 0 36 0 0 110 4
1789 1111
1789 1072
1645 1072
1645 532
3 2 12 0 0 12416 0 36 0 0 110 4
1834 1111
1834 1067
1655 1067
1655 532
1 8 13 0 0 4224 0 0 35 110 0 4
2047 532
2047 1067
1927 1067
1927 1111
3 0 14 0 0 12416 0 35 0 0 110 4
1972 1111
1972 1073
2061 1073
2061 532
8 7 15 0 0 4096 0 33 0 0 110 2
1789 810
1789 532
3 6 16 0 0 4096 0 33 0 0 110 2
1834 810
1834 532
8 5 17 0 0 4096 0 34 0 0 110 2
1928 810
1928 532
3 4 18 0 0 4096 0 34 0 0 110 2
1973 810
1973 532
16 7 15 0 0 0 0 72 0 0 110 2
364 510
364 532
15 6 16 0 0 0 0 72 0 0 110 2
373 510
373 532
14 5 17 0 0 0 0 72 0 0 110 2
382 510
382 532
13 4 18 0 0 0 0 72 0 0 110 2
391 510
391 532
12 3 11 0 0 0 0 72 0 0 110 2
409 510
409 532
11 2 12 0 0 0 0 72 0 0 110 2
418 510
418 532
10 1 13 0 0 0 0 72 0 0 110 2
427 510
427 532
9 0 14 0 0 0 0 72 0 0 110 2
436 510
436 532
1 1 19 0 0 12416 0 72 42 0 0 4
436 446
436 431
463 431
463 400
2 2 20 0 0 8320 0 72 42 0 0 4
427 446
427 426
457 426
457 400
3 3 21 0 0 8320 0 72 42 0 0 4
418 446
418 421
451 421
451 400
4 4 22 0 0 8320 0 72 42 0 0 4
409 446
409 417
445 417
445 400
4 8 23 0 0 4224 0 20 72 0 0 2
364 401
364 446
3 7 24 0 0 4224 0 20 72 0 0 4
370 401
370 426
373 426
373 446
2 6 25 0 0 12416 0 20 72 0 0 4
376 401
376 421
382 421
382 446
5 1 26 0 0 4224 0 72 20 0 0 4
391 446
391 417
382 417
382 401
1 1 27 0 0 12416 0 5 71 0 0 4
314 759
334 759
334 758
404 758
1 2 2 0 0 0 0 70 5 0 0 3
273 787
273 759
280 759
3 1 8 0 0 0 0 71 2 0 0 6
455 767
501 767
501 808
387 808
387 854
404 854
4 2 28 0 0 12416 0 2 71 0 0 6
455 863
503 863
503 820
394 820
394 776
404 776
1 1 4 0 0 0 3 14 6 0 0 3
1221 362
1221 363
1510 363
0 1 29 0 0 8192 0 0 10 46 0 4
987 229
987 230
1495 230
1495 261
0 1 29 0 0 4224 0 0 13 121 0 5
796 748
796 229
989 229
989 261
990 261
6 1 30 0 0 12416 0 9 18 0 0 5
1750 389
1761 389
1761 504
704 504
704 407
2 6 31 0 0 8320 0 18 8 0 0 5
698 407
698 511
1687 511
1687 389
1677 389
6 3 32 0 0 12416 0 7 18 0 0 5
1607 389
1616 389
1616 517
692 517
692 407
4 6 33 0 0 8320 0 18 6 0 0 5
686 407
686 524
1546 524
1546 390
1534 390
6 1 34 0 0 12416 0 14 19 0 0 7
1245 389
1258 389
1258 469
641 469
641 417
619 417
619 408
2 6 35 0 0 16512 0 19 15 0 0 9
613 408
613 423
634 423
634 475
1183 475
1183 388
1176 388
1176 389
1172 389
3 6 36 0 0 16512 0 19 16 0 0 7
607 408
607 427
630 427
630 481
1111 481
1111 389
1102 389
6 4 37 0 0 12416 0 17 19 0 0 5
1029 390
1040 390
1040 491
601 491
601 408
2 4 18 0 0 12288 0 13 0 0 110 4
981 261
981 221
843 221
843 532
4 5 17 0 0 12288 0 13 0 0 110 4
963 261
963 216
833 216
833 532
6 6 16 0 0 12288 0 13 0 0 110 4
945 261
945 212
823 212
823 532
8 7 15 0 0 12288 0 13 0 0 110 4
927 261
927 209
814 209
814 532
2 0 14 0 0 0 0 10 0 0 110 4
1486 261
1486 222
1379 222
1379 532
4 1 13 0 0 0 0 10 0 0 110 4
1468 261
1468 215
1373 215
1373 532
6 2 12 0 0 0 0 10 0 0 110 4
1450 261
1450 208
1367 208
1367 532
8 3 11 0 0 0 0 10 0 0 110 4
1432 261
1432 203
1363 203
1363 532
0 4 4 0 0 0 0 0 6 70 0 2
1510 443
1510 438
3 0 38 0 0 8192 0 7 0 0 65 3
1559 407
1550 407
1550 454
0 0 38 0 0 4096 0 0 0 67 66 4
1622 454
1451 454
1451 453
1447 453
3 0 38 0 0 12288 0 6 0 0 84 4
1486 408
1447 408
1447 454
1187 454
3 3 38 0 0 0 0 8 9 0 0 6
1629 407
1622 407
1622 454
1692 454
1692 407
1702 407
0 4 4 0 0 0 0 0 9 69 0 3
1652 443
1726 443
1726 437
0 4 4 0 0 0 0 0 8 70 0 3
1583 443
1653 443
1653 437
0 4 4 0 0 0 0 0 7 86 0 3
1221 443
1583 443
1583 437
1 1 4 0 0 0 3 8 9 0 0 4
1653 362
1653 363
1726 363
1726 362
1 1 4 0 0 0 3 7 8 0 0 4
1583 362
1583 363
1653 363
1653 362
1 1 4 0 0 0 3 6 7 0 0 3
1510 363
1583 363
1583 362
6 3 30 0 0 0 0 9 10 0 0 4
1750 389
1750 242
1477 242
1477 261
6 5 31 0 0 0 0 8 10 0 0 4
1677 389
1677 247
1459 247
1459 261
6 7 32 0 0 0 0 7 10 0 0 4
1607 389
1607 251
1441 251
1441 261
6 9 33 0 0 0 0 6 10 0 0 4
1534 390
1534 255
1423 255
1423 261
1 10 2 0 0 0 0 11 10 0 0 4
1414 255
1414 252
1414 252
1414 255
11 2 39 0 0 8320 0 10 9 0 0 5
1477 325
1477 328
1692 328
1692 389
1702 389
12 2 40 0 0 8320 0 10 8 0 0 5
1459 325
1459 333
1621 333
1621 389
1629 389
13 2 41 0 0 8320 0 10 7 0 0 5
1441 325
1441 339
1550 339
1550 389
1559 389
14 2 42 0 0 4224 0 10 6 0 0 3
1423 325
1423 390
1486 390
3 0 38 0 0 0 0 17 0 0 85 3
981 408
946 408
946 454
0 3 38 0 0 0 0 0 14 85 0 4
1116 454
1187 454
1187 407
1197 407
0 3 38 0 0 4096 0 0 15 164 0 5
601 1282
601 454
1116 454
1116 407
1124 407
0 4 4 0 0 0 0 0 14 87 0 3
1147 443
1221 443
1221 437
0 4 4 0 0 0 0 0 15 88 0 3
1078 443
1148 443
1148 437
0 4 4 0 0 0 0 0 16 128 0 3
1005 443
1078 443
1078 437
1 1 4 0 0 0 3 15 14 0 0 4
1148 362
1148 363
1221 363
1221 362
1 1 4 0 0 0 3 16 15 0 0 4
1078 362
1078 363
1148 363
1148 362
1 1 4 0 0 0 3 17 16 0 0 3
1005 363
1078 363
1078 362
0 1 4 0 0 4096 3 0 17 178 0 5
589 1020
589 673
787 673
787 363
1005 363
6 3 34 0 0 0 0 14 13 0 0 4
1245 389
1245 242
972 242
972 261
6 5 35 0 0 0 0 15 13 0 0 4
1172 389
1172 247
954 247
954 261
6 7 36 0 0 0 0 16 13 0 0 4
1102 389
1102 251
936 251
936 261
6 9 37 0 0 0 0 17 13 0 0 4
1029 390
1029 255
918 255
918 261
1 10 2 0 0 0 0 12 13 0 0 4
909 255
909 252
909 252
909 255
11 2 43 0 0 8320 0 13 14 0 0 5
972 325
972 328
1187 328
1187 389
1197 389
12 2 44 0 0 8320 0 13 15 0 0 5
954 325
954 333
1116 333
1116 389
1124 389
13 2 45 0 0 8320 0 13 16 0 0 5
936 325
936 339
1045 339
1045 389
1054 389
14 2 46 0 0 4224 0 13 17 0 0 3
918 325
918 390
981 390
9 7 15 0 0 8320 0 69 0 0 110 3
2314 868
2318 868
2318 532
10 6 16 0 0 8320 0 69 0 0 110 3
2314 877
2326 877
2326 532
11 5 17 0 0 8320 0 69 0 0 110 3
2314 886
2338 886
2338 532
12 4 18 0 0 8320 0 69 0 0 110 3
2314 895
2345 895
2345 532
13 3 11 0 0 0 0 69 0 0 110 3
2314 913
2354 913
2354 532
14 2 12 0 0 0 0 69 0 0 110 3
2314 922
2365 922
2365 532
1 15 13 0 0 0 0 0 69 110 0 3
2375 532
2375 931
2314 931
16 0 14 0 0 0 0 69 0 0 110 3
2314 940
2386 940
2386 532
-215140 0 1 0 0 4256 0 0 0 0 0 2
272 532
2554 532
17 0 47 0 0 4096 0 69 0 0 112 2
2244 859
2224 859
5 18 47 0 0 12416 0 68 69 0 0 6
896 1153
962 1153
962 695
2224 695
2224 904
2244 904
0 5 48 0 0 4224 0 0 69 240 0 4
1796 885
2182 885
2182 913
2250 913
0 6 49 0 0 4224 0 0 69 238 0 4
1870 889
2175 889
2175 922
2250 922
0 7 50 0 0 4224 0 0 69 236 0 4
1940 895
2170 895
2170 931
2250 931
8 0 51 0 0 4224 0 69 0 0 261 2
2250 940
2095 940
1 0 2 0 0 0 0 69 0 0 119 2
2250 868
2238 868
2 0 2 0 0 0 0 69 0 0 119 2
2250 877
2238 877
0 3 2 0 0 4224 0 0 69 241 0 4
1955 789
2238 789
2238 886
2250 886
0 4 52 0 0 4096 0 0 69 253 0 3
2193 1087
2193 895
2250 895
6 1 29 0 0 0 0 68 57 0 0 6
890 1135
942 1135
942 748
785 748
785 799
791 799
1 0 53 0 0 4096 0 47 0 0 167 3
756 1126
702 1126
702 1104
1 2 54 0 0 8192 0 45 47 0 0 4
670 722
681 722
681 1144
756 1144
3 2 55 0 0 4224 0 47 68 0 0 2
801 1135
842 1135
3 0 56 0 0 4096 0 68 0 0 175 2
842 1153
828 1153
1 0 4 0 0 0 3 68 0 0 161 2
866 1108
610 1108
4 0 4 0 0 0 0 53 0 0 128 2
866 1096
950 1096
0 4 4 0 0 12416 0 0 17 179 0 6
950 982
950 1253
617 1253
617 443
1005 443
1005 438
1 0 53 0 0 0 0 67 0 0 131 3
2453 1209
2454 1209
2454 1197
2 2 57 0 0 4224 0 65 67 0 0 3
2437 1259
2453 1259
2453 1245
0 1 53 0 0 4224 0 0 64 194 0 4
1548 999
2454 999
2454 1197
2440 1197
3 2 58 0 0 4224 0 28 64 0 0 4
2338 1151
2445 1151
2445 1179
2440 1179
0 1 52 0 0 8320 0 0 65 254 0 5
2191 1227
2191 1299
2451 1299
2451 1277
2437 1277
3 2 59 0 0 4224 0 66 31 0 0 2
2334 1227
2290 1227
1 3 60 0 0 8320 0 66 65 0 0 3
2380 1236
2392 1236
2392 1268
3 2 61 0 0 4224 0 64 66 0 0 3
2395 1188
2395 1218
2380 1218
1 1 4 0 0 0 3 59 32 0 0 2
1436 899
1353 899
2 5 62 0 0 4224 0 58 59 0 0 4
1243 713
1482 713
1482 944
1466 944
6 1 63 0 0 8320 0 43 58 0 0 4
1290 927
1307 927
1307 731
1243 731
3 0 64 0 0 4096 0 59 0 0 188 3
1412 944
1412 1061
1329 1061
0 4 4 0 0 0 0 0 59 189 0 3
1353 981
1436 981
1436 974
3 2 65 0 0 8320 0 63 59 0 0 4
1418 1002
1402 1002
1402 926
1412 926
1 0 66 0 0 8320 0 63 0 0 146 4
1463 1011
1463 1053
1270 1053
1270 1035
5 2 62 0 0 0 0 59 63 0 0 3
1466 944
1466 993
1463 993
3 2 67 0 0 4224 0 62 32 0 0 3
1311 986
1311 926
1329 926
0 1 66 0 0 0 0 0 62 152 0 4
1270 999
1270 1035
1302 1035
1302 1031
3 2 68 0 0 4224 0 61 62 0 0 3
1354 1034
1320 1034
1320 1031
0 2 69 0 0 8192 0 0 61 151 0 4
1394 926
1406 926
1406 1025
1403 1025
0 1 70 0 0 4096 0 0 61 150 0 3
1475 926
1475 1043
1403 1043
6 1 70 0 0 12416 0 59 60 0 0 5
1460 926
1475 926
1475 893
1174 893
1174 918
2 6 69 0 0 12416 0 60 32 0 0 6
1174 927
1168 927
1168 888
1394 888
1394 926
1377 926
5 3 66 0 0 0 0 43 60 0 0 5
1296 945
1296 999
1168 999
1168 936
1174 936
4 2 71 0 0 4224 0 60 43 0 0 2
1219 927
1242 927
0 7 72 0 0 8192 0 0 35 211 0 4
1871 1101
1871 1084
1936 1084
1936 1111
7 0 2 0 0 0 0 36 0 0 216 2
1798 1111
1798 1090
0 0 7 0 0 4224 0 0 0 197 170 4
1636 805
994 805
994 926
928 926
4 0 4 0 0 0 0 43 0 0 189 2
1266 975
1266 981
1 3 54 0 0 4224 0 45 58 0 0 2
670 722
1198 722
0 0 53 0 0 0 0 0 0 195 194 2
1762 798
1548 798
12 0 7 0 0 0 0 33 0 0 197 2
1753 810
1753 805
0 0 4 0 0 8320 3 0 0 178 249 3
610 1020
610 1198
1575 1198
4 4 4 0 0 0 0 21 22 0 0 4
1772 966
1772 977
1846 977
1846 972
4 0 4 0 0 0 0 21 0 0 203 4
1772 966
1772 976
1599 976
1599 1278
4 0 38 0 0 16512 0 49 0 0 202 5
340 1200
340 1282
621 1282
621 1283
1667 1283
3 0 38 0 0 0 0 41 0 0 202 3
1749 1244
1737 1244
1737 1283
0 3 64 0 0 4224 0 0 48 188 0 2
1242 1061
1060 1061
2 0 53 0 0 0 0 44 0 0 174 5
690 1076
626 1076
626 1104
924 1104
924 1048
1 2 73 0 0 8320 0 44 45 0 0 4
690 1058
627 1058
627 722
634 722
2 3 74 0 0 4224 0 46 44 0 0 4
774 1057
745 1057
745 1067
735 1067
6 1 7 0 0 0 0 52 46 0 0 6
887 926
928 926
928 990
728 990
728 1039
774 1039
3 2 75 0 0 4224 0 46 53 0 0 2
820 1048
842 1048
1 1 4 0 0 0 3 52 43 0 0 4
863 899
863 898
1266 898
1266 900
0 2 56 0 0 4096 0 0 48 175 0 4
828 1191
1002 1191
1002 1070
1015 1070
1 6 53 0 0 0 0 48 53 0 0 4
1015 1052
1003 1052
1003 1048
890 1048
3 0 56 0 0 4224 0 49 0 0 181 5
334 1191
828 1191
828 1107
830 1107
830 1065
4 0 4 0 0 0 3 51 0 0 177 3
863 856
808 856
808 898
1 0 4 0 0 0 3 52 0 0 178 4
863 899
863 898
808 898
808 1020
1 1 4 0 0 0 3 50 53 0 0 7
279 1020
428 1020
428 1019
589 1019
589 1020
866 1020
866 1021
4 1 4 0 0 0 0 52 51 0 0 6
863 974
863 982
950 982
950 759
863 759
863 781
3 0 56 0 0 0 0 52 0 0 181 2
839 944
830 944
3 3 56 0 0 0 0 53 51 0 0 5
842 1066
842 1065
830 1065
830 826
839 826
3 2 76 0 0 4224 0 54 57 0 0 3
792 816
792 817
791 817
3 2 77 0 0 4224 0 57 51 0 0 4
837 808
840 808
840 808
839 808
2 0 78 0 0 8192 0 54 0 0 186 4
747 825
737 825
737 888
736 888
2 1 79 0 0 4224 0 56 54 0 0 2
727 807
747 807
6 1 78 0 0 12416 0 51 55 0 0 6
887 808
935 808
935 888
736 888
736 917
749 917
3 2 80 0 0 4224 0 55 52 0 0 2
794 926
839 926
3 3 64 0 0 0 0 32 43 0 0 4
1329 944
1329 1061
1242 1061
1242 945
0 4 4 0 0 0 0 0 32 128 0 5
950 1179
1159 1179
1159 981
1353 981
1353 974
1 1 4 0 0 0 3 43 32 0 0 4
1266 900
1266 898
1353 898
1353 899
3 7 81 0 0 8320 0 29 33 0 0 4
2332 1078
2332 785
1798 785
1798 810
0 1 72 0 0 0 0 0 36 211 0 2
1852 1101
1852 1111
11 11 53 0 0 0 0 36 35 0 0 4
1762 1111
1762 1096
1900 1096
1900 1111
11 0 53 0 0 0 0 36 0 0 174 6
1762 1111
1762 1096
1548 1096
1548 797
972 797
972 1048
11 11 53 0 0 0 0 33 34 0 0 4
1762 810
1762 797
1901 797
1901 810
12 12 7 0 0 0 0 36 35 0 0 4
1753 1111
1753 1107
1891 1107
1891 1111
12 12 7 0 0 0 0 36 34 0 0 6
1753 1111
1753 1107
1636 1107
1636 805
1892 805
1892 810
2 0 82 0 0 12288 0 26 0 0 208 4
2141 1078
2094 1078
2094 1101
2020 1101
1 1 4 0 0 0 3 31 38 0 0 3
2266 1200
2266 1198
1989 1198
0 3 38 0 0 0 0 0 31 223 0 4
1959 1284
2328 1284
2328 1245
2290 1245
3 0 38 0 0 0 0 22 0 0 252 3
1822 942
1814 942
1814 983
3 3 38 0 0 0 0 21 40 0 0 6
1748 936
1667 936
1667 1283
1816 1283
1816 1243
1822 1243
0 0 4 0 0 0 0 0 0 189 204 3
1159 1178
1159 1278
1773 1278
4 4 4 0 0 0 0 41 40 0 0 4
1773 1274
1773 1278
1846 1278
1846 1273
2 0 83 0 0 8192 0 35 0 0 209 3
1981 1111
1981 1105
1946 1105
0 2 84 0 0 4096 0 0 36 212 0 3
1807 1104
1843 1104
1843 1111
0 4 82 0 0 0 0 0 35 208 0 3
1991 1101
1963 1101
1963 1111
6 1 82 0 0 8320 0 38 35 0 0 5
2013 1225
2020 1225
2020 1101
1990 1101
1990 1111
0 6 83 0 0 0 0 0 35 210 0 5
1919 1101
1946 1101
1946 1105
1945 1105
1945 1111
6 9 83 0 0 16512 0 39 35 0 0 9
1940 1225
1941 1225
1941 1177
1877 1177
1877 1101
1919 1101
1919 1101
1918 1101
1918 1111
6 4 72 0 0 8320 0 40 36 0 0 5
1870 1225
1871 1225
1871 1101
1825 1101
1825 1111
0 6 84 0 0 0 0 0 36 213 0 3
1779 1101
1807 1101
1807 1111
6 9 84 0 0 12416 0 41 36 0 0 6
1797 1226
1797 1179
1735 1179
1735 1101
1780 1101
1780 1111
5 0 2 0 0 0 0 35 0 0 215 3
1954 1105
1954 1090
1910 1090
10 0 2 0 0 0 0 35 0 0 216 5
1909 1105
1909 1090
1910 1090
1910 1090
1816 1090
5 0 2 0 0 0 0 36 0 0 217 3
1816 1105
1816 1090
1771 1090
10 1 2 0 0 0 0 36 37 0 0 3
1771 1105
1771 1090
1735 1090
14 2 85 0 0 12416 0 35 38 0 0 5
1972 1175
1972 1184
1953 1184
1953 1225
1965 1225
13 2 86 0 0 8320 0 35 39 0 0 5
1927 1175
1927 1184
1884 1184
1884 1225
1892 1225
14 2 87 0 0 12416 0 36 40 0 0 5
1834 1175
1834 1186
1815 1186
1815 1225
1822 1225
13 2 88 0 0 8320 0 36 41 0 0 5
1789 1175
1789 1184
1737 1184
1737 1226
1749 1226
4 0 4 0 0 0 0 41 0 0 204 2
1773 1274
1773 1278
0 3 38 0 0 0 0 0 38 224 0 4
1888 1284
1959 1284
1959 1243
1965 1243
0 3 38 0 0 0 0 0 39 202 0 6
1816 1283
1822 1283
1822 1284
1888 1284
1888 1243
1892 1243
0 4 4 0 0 0 0 0 38 226 0 3
1915 1279
1989 1279
1989 1273
0 4 4 0 0 0 0 0 39 204 0 4
1846 1278
1846 1279
1916 1279
1916 1273
1 1 4 0 0 0 3 39 38 0 0 2
1916 1198
1989 1198
1 1 4 0 0 0 3 40 39 0 0 2
1846 1198
1916 1198
1 1 4 0 0 0 3 41 40 0 0 3
1773 1199
1773 1198
1846 1198
2 0 50 0 0 0 0 34 0 0 235 3
1982 810
1982 804
1946 804
7 0 49 0 0 0 0 34 0 0 238 3
1937 810
1937 802
1870 802
0 2 48 0 0 0 0 0 33 239 0 3
1807 803
1843 803
1843 810
0 4 51 0 0 0 0 0 34 234 0 3
1991 800
1964 800
1964 810
0 1 51 0 0 0 0 0 34 261 0 4
2019 924
2019 800
1991 800
1991 810
0 6 50 0 0 0 0 0 34 236 0 3
1919 800
1946 800
1946 810
6 9 50 0 0 0 0 23 34 0 0 6
1940 924
1940 878
1880 878
1880 800
1919 800
1919 810
0 4 49 0 0 0 0 0 33 238 0 3
1852 800
1825 800
1825 810
6 1 49 0 0 0 0 22 33 0 0 4
1870 924
1870 800
1852 800
1852 810
0 6 48 0 0 0 0 0 33 240 0 3
1779 800
1807 800
1807 810
6 9 48 0 0 0 0 21 33 0 0 8
1796 918
1796 880
1797 880
1797 878
1735 878
1735 800
1780 800
1780 810
5 0 2 0 0 0 0 34 0 0 242 3
1955 804
1955 789
1910 789
10 0 2 0 0 0 0 34 0 0 243 3
1910 804
1910 789
1816 789
5 0 2 0 0 0 0 33 0 0 244 3
1816 804
1816 789
1771 789
10 1 2 0 0 0 0 33 25 0 0 3
1771 804
1771 789
1735 789
14 2 89 0 0 12416 0 34 24 0 0 5
1973 874
1973 883
1953 883
1953 924
1965 924
13 2 90 0 0 8320 0 34 23 0 0 5
1928 874
1928 883
1884 883
1884 924
1892 924
14 2 91 0 0 12416 0 33 22 0 0 5
1834 874
1834 885
1815 885
1815 924
1822 924
13 2 92 0 0 8320 0 33 21 0 0 5
1789 874
1789 883
1737 883
1737 918
1748 918
1 1 4 0 0 0 3 21 41 0 0 5
1772 891
1575 891
1575 1198
1773 1198
1773 1199
4 0 4 0 0 0 0 21 0 0 162 4
1772 966
1772 975
1773 975
1773 977
0 3 38 0 0 0 0 0 24 252 0 4
1892 983
1959 983
1959 942
1965 942
0 3 38 0 0 0 0 0 23 202 0 3
1667 983
1892 983
1892 942
2 0 52 0 0 0 0 29 0 0 254 3
2283 1087
2191 1087
2191 1184
6 2 52 0 0 0 0 31 30 0 0 4
2242 1227
2191 1227
2191 1184
2221 1184
1 0 93 0 0 8320 0 30 0 0 258 3
2221 1166
2210 1166
2210 1069
2 3 94 0 0 8320 0 28 30 0 0 4
2287 1160
2282 1160
2282 1175
2272 1175
3 1 95 0 0 8320 0 27 28 0 0 4
2271 1128
2281 1128
2281 1142
2287 1142
3 1 93 0 0 0 0 26 29 0 0 2
2190 1069
2283 1069
2 0 82 0 0 0 0 27 0 0 198 3
2220 1137
2134 1137
2134 1078
0 1 51 0 0 0 0 0 27 261 0 3
2123 1060
2123 1119
2220 1119
6 1 51 0 0 0 0 24 26 0 0 4
2013 924
2095 924
2095 1060
2141 1060
0 4 4 0 0 0 0 0 24 263 0 3
1915 978
1989 978
1989 972
0 4 4 0 0 0 0 0 23 162 0 4
1846 977
1846 978
1916 978
1916 972
1 1 4 0 0 0 3 23 24 0 0 4
1916 897
1916 898
1989 898
1989 897
1 1 4 0 0 0 3 22 23 0 0 4
1846 897
1846 898
1916 898
1916 897
1 1 4 0 0 0 3 21 22 0 0 4
1772 891
1772 892
1846 892
1846 897
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2320 1046 2391 1070
2340 1062 2370 1078
3 SUM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2072 1156 2203 1180
2092 1172 2182 1188
9 CARRY BIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2320 1090 2461 1114
2340 1106 2440 1122
10 FULL ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
576 282 727 306
596 298 706 314
11 OUTPUT UNIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1180 98 1341 122
1200 114 1320 130
12 SERIAL ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1512 213 1619 237
1517 217 1613 233
12 REGISTER LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
971 194 1066 218
982 202 1054 218
12 REGISTER MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
691 1216 806 1237
700 1222 796 1237
12 CONTROL UNIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1576 759 1635 781
1585 766 1625 782
5 SHIFT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1576 811 1627 833
1585 819 1617 835
4 LOAD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1828 728 1927 743
1842 740 1912 751
10 REGISTER A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1829 1040 1930 1055
1844 1051 1914 1062
10 REGISTER B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
1142 849 1281 871
1151 856 1271 872
15 MOD - 5 COUNTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
367 297 466 319
376 304 456 320
10 INPUT UNIT
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
