CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 60 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
67
8 SPDT PB~
217 150 426 0 10 18
0 7 3 2 0 0 0 0 0 0
1
0
0 0 4704 0
0
5 RESET
-14 -15 21 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
5130 0 0
2
5.89984e-315 0
0
5 7474~
219 1055 760 0 6 22
0 3 95 4 7 96 87
0
0 0 4704 0
4 7474
7 -60 35 -52
2 R7
-8 -31 6 -23
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
391 0 0
2
44326.5 0
0
5 7474~
219 1129 760 0 6 22
0 3 94 4 7 97 86
0
0 0 4704 0
4 7474
7 -60 35 -52
2 R6
-6 -33 8 -25
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
3124 0 0
2
44326.5 1
0
5 7474~
219 1199 760 0 6 22
0 3 93 4 7 98 85
0
0 0 4704 0
4 7474
7 -60 35 -52
2 R5
-7 -32 7 -24
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
3421 0 0
2
44326.5 2
0
5 7474~
219 1271 760 0 6 22
0 3 92 4 7 99 84
0
0 0 4704 0
4 7474
7 -60 35 -52
2 R4
-7 -32 7 -24
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
8157 0 0
2
44326.5 3
0
7 Ground~
168 973 567 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
44326.5 4
0
4 4539
219 1091 636 0 14 29
0 86 63 87 86 2 87 64 2 87
2 41 12 95 94
0
0 0 4320 270
4 4539
-14 -60 14 -52
3 U17
62 9 83 17
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
8901 0 0
2
44326.5 5
0
4 4539
219 1230 636 0 14 29
0 84 61 85 84 2 85 62 86 85
2 41 12 93 92
0
0 0 4320 270
4 4539
-14 -60 14 -52
3 U13
62 9 83 17
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
7361 0 0
2
44326.5 6
0
4 4539
219 1515 635 0 14 29
0 44 57 81 44 2 81 58 82 81
2 41 12 89 88
0
0 0 4320 270
4 4539
-14 -60 14 -52
2 U3
65 9 79 17
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
44326.5 7
0
4 4539
219 1376 635 0 14 29
0 82 59 83 82 2 83 60 84 83
2 41 12 91 90
0
0 0 4320 270
4 4539
-14 -60 14 -52
2 U4
65 9 79 17
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
44326.5 8
0
5 7474~
219 1557 760 0 6 22
0 3 88 4 7 100 44
0
0 0 4704 0
4 7474
7 -60 35 -52
2 R0
-8 -31 6 -23
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
3472 0 0
2
44326.5 9
0
5 7474~
219 1484 760 0 6 22
0 3 89 4 7 101 81
0
0 0 4704 0
4 7474
7 -60 35 -52
2 R1
-6 -32 8 -24
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 3 0
1 U
9998 0 0
2
44326.5 10
0
5 7474~
219 1414 760 0 6 22
0 3 90 4 7 102 82
0
0 0 4704 0
4 7474
7 -60 35 -52
2 R2
-7 -32 7 -24
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
3536 0 0
2
44326.5 11
0
5 7474~
219 1340 760 0 6 22
0 3 91 4 7 103 83
0
0 0 4704 0
4 7474
7 -60 35 -52
2 R3
-6 -32 8 -24
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 4 0
1 U
4597 0 0
2
44326.5 12
0
5 7474~
219 548 526 0 6 22
0 7 77 15 3 104 74
0
0 0 4704 0
4 7474
7 -60 35 -52
2 T1
-8 -31 6 -23
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 5 0
1 U
3835 0 0
2
44326.5 13
0
5 7474~
219 548 626 0 6 22
0 3 73 15 7 6 41
0
0 0 4704 0
4 7474
7 -60 35 -52
2 T2
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 5 0
1 U
3670 0 0
2
44326.5 14
0
5 7474~
219 546 732 0 6 22
0 3 42 15 7 105 29
0
0 0 4704 0
4 7474
7 -60 35 -52
2 T3
-7 -31 7 -23
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 6 0
1 U
5616 0 0
2
44326.5 15
0
5 7474~
219 545 835 0 6 22
0 3 38 15 7 106 12
0
0 0 4704 0
4 7474
7 -60 35 -52
2 T4
-7 -32 7 -24
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 6 0
1 U
9323 0 0
2
44326.5 16
0
5 7474~
219 544 937 0 6 22
0 3 37 15 7 107 16
0
0 0 4704 0
4 7474
7 -60 35 -52
2 T5
-6 -33 8 -25
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 7 0
1 U
317 0 0
2
44326.5 17
0
5 7474~
219 544 1039 0 6 22
0 3 34 15 7 25 24
0
0 0 4704 0
4 7474
7 -60 35 -52
2 T6
-6 -32 8 -24
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 7 0
1 U
3108 0 0
2
44326.5 18
0
14 NO PushButton~
191 152 473 0 2 5
0 80 2
0
0 0 4704 0
0
5 COUNT
-17 -20 18 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4299 0 0
2
44326.5 19
0
10 2-In NAND~
219 266 490 0 3 22
0 80 79 75
0
0 0 96 0
6 74LS00
-14 -24 28 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
9672 0 0
2
44326.5 20
0
7 Ground~
168 91 518 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7876 0 0
2
44326.5 21
0
5 4023~
219 267 560 0 4 22
0 75 7 6 79
0
0 0 96 0
4 4023
-14 -28 14 -20
4 U11A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 9 0
1 U
6369 0 0
2
44326.5 22
0
8 2-In OR~
219 460 490 0 3 22
0 24 78 77
0
0 0 96 0
6 74LS32
-21 -24 21 -16
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
9172 0 0
2
44326.5 23
0
9 2-In AND~
219 399 499 0 3 22
0 76 74 78
0
0 0 96 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
7100 0 0
2
44326.5 24
0
9 2-In AND~
219 471 590 0 3 22
0 74 75 73
0
0 0 96 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3820 0 0
2
44326.5 25
0
9 Inverter~
13 348 490 0 2 22
0 75 76
0
0 0 96 0
6 74LS04
-21 -19 21 -11
4 U15A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
7678 0 0
2
44326.5 26
0
2 +V
167 92 555 0 1 3
0 3
0
0 0 54112 0
2 5V
-7 -14 7 -6
3 VCC
-10 -24 11 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
961 0 0
2
44326.5 27
0
8 Hex Key~
166 169 276 0 11 12
0 69 70 71 72 0 0 0 0 0
0 48
0
0 0 4640 0
0
3 MSB
-11 -34 10 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3178 0 0
2
44326.5 28
0
8 Hex Key~
166 215 275 0 11 12
0 65 66 67 68 0 0 0 0 0
0 48
0
0 0 4640 0
0
3 LSB
-11 -34 10 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3409 0 0
2
44326.5 29
0
7 74LS244
143 202 341 0 18 37
0 65 66 67 68 69 70 71 72 57
58 59 60 61 62 63 64 6 6
0
0 0 4320 270
6 74F244
-21 -60 21 -52
2 U2
54 0 68 8
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 0 0 0
1 U
3951 0 0
2
44326.5 30
0
7 Ground~
168 430 141 0 1 3
0 2
0
0 0 53344 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8885 0 0
2
44326.5 31
0
7 74LS157
122 476 182 0 14 29
0 24 23 52 22 51 21 50 20 49
2 53 54 55 56
0
0 0 4320 270
6 74F157
-21 -60 21 -52
3 U24
51 0 72 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3780 0 0
2
44326.5 32
0
5 7474~
219 742 319 0 6 22
0 3 53 4 7 108 52
0
0 0 4192 0
4 7474
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 13 0
1 U
9265 0 0
2
44326.5 33
0
5 7474~
219 669 319 0 6 22
0 3 54 4 7 109 51
0
0 0 4192 0
4 7474
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 13 0
1 U
9442 0 0
2
44326.5 34
0
5 7474~
219 599 319 0 6 22
0 3 55 4 7 110 50
0
0 0 4192 0
4 7474
7 -60 35 -52
3 U5A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 14 0
1 U
9424 0 0
2
44326.5 35
0
5 7474~
219 526 320 0 6 22
0 3 56 4 7 111 49
0
0 0 4192 0
4 7474
7 -60 35 -52
3 U5B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 14 0
1 U
9968 0 0
2
44326.5 36
0
12 Hex Display~
7 390 276 0 16 19
10 52 51 50 49 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 COUNT
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9281 0 0
2
44326.5 37
0
9 2-In AND~
219 1417 874 0 3 22
0 44 29 48
0
0 0 96 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
8464 0 0
2
44326.5 38
0
9 2-In AND~
219 1417 937 0 3 22
0 45 43 47
0
0 0 96 0
6 74LS08
-21 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
7168 0 0
2
44326.5 39
0
5 7474~
219 1555 942 0 6 22
0 3 46 4 7 35 43
0
0 0 4704 0
4 7474
7 -60 35 -52
4 FLAG
-14 -31 14 -23
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 15 0
1 U
3171 0 0
2
44326.5 40
0
8 2-In OR~
219 1479 905 0 3 22
0 48 47 46
0
0 0 96 0
6 74LS32
-21 -24 21 -16
4 U12B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
4139 0 0
2
44326.5 41
0
9 Inverter~
13 1308 928 0 2 22
0 29 45
0
0 0 96 0
6 74LS04
-21 -19 21 -11
4 U15B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
6435 0 0
2
44326.5 42
0
8 3-In OR~
219 455 696 0 4 22
0 41 40 39 42
0
0 0 96 0
4 4075
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 18 0
1 U
5283 0 0
2
44326.5 43
0
9 2-In AND~
219 401 696 0 3 22
0 35 12 40
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 19 0
1 U
6874 0 0
2
44326.5 44
0
9 2-In AND~
219 400 734 0 3 22
0 16 31 39
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 19 0
1 U
5305 0 0
2
44326.5 45
0
9 2-In AND~
219 469 799 0 3 22
0 31 29 38
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
34 0 0
2
44326.5 46
0
9 2-In AND~
219 468 901 0 3 22
0 12 36 37
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
969 0 0
2
44326.5 47
0
9 Inverter~
13 404 911 0 2 22
0 35 36
0
0 0 96 0
6 74LS04
-21 -19 21 -11
4 U15C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 12 0
1 U
8402 0 0
2
44326.5 48
0
8 2-In OR~
219 457 1003 0 3 22
0 33 32 34
0
0 0 96 0
6 74LS32
-21 -24 21 -16
4 U12C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
3751 0 0
2
44326.5 49
0
9 2-In AND~
219 403 979 0 3 22
0 29 30 33
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
4292 0 0
2
44326.5 50
0
9 2-In AND~
219 405 1027 0 3 22
0 30 16 32
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 20 0
1 U
6118 0 0
2
44326.5 51
0
9 Inverter~
13 647 826 0 2 22
0 31 30
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 U15D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
34 0 0
2
44326.5 52
0
7 74LS125
115 1887 591 0 12 25
0 25 28 25 17 25 27 25 26 23
22 21 20
0
0 0 4320 90
6 74F125
-21 -51 21 -43
2 U9
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
6357 0 0
2
44326.5 53
0
6 74112~
219 717 918 0 7 32
0 3 12 15 12 5 19 11
0
0 0 4704 0
5 74112
4 -60 39 -52
2 Q0
-8 -22 6 -14
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 16 0
1 U
319 0 0
2
44326.5 54
0
6 74112~
219 802 920 0 7 32
0 3 12 19 12 5 18 10
0
0 0 4704 0
5 74112
4 -60 39 -52
2 Q1
-9 -19 5 -11
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 16 0
1 U
3976 0 0
2
44326.5 55
0
6 74112~
219 883 917 0 7 32
0 3 12 18 12 5 13 9
0
0 0 4704 0
5 74112
4 -60 39 -52
2 Q2
-7 -22 7 -14
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 16 0
1 U
7634 0 0
2
44326.5 56
0
6 74112~
219 1749 760 0 7 32
0 3 16 15 16 14 112 28
0
0 0 4704 0
5 74112
4 -60 39 -52
2 Q0
-6 -20 8 -12
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 17 0
1 U
523 0 0
2
44326.5 57
0
6 74112~
219 1827 759 0 7 32
0 3 16 28 16 14 113 17
0
0 0 4704 0
5 74112
4 -60 39 -52
2 Q1
-6 -20 8 -12
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 17 0
1 U
6748 0 0
2
44326.5 58
0
6 74112~
219 1899 759 0 7 32
0 3 16 17 16 14 114 27
0
0 0 4704 0
5 74112
4 -60 39 -52
2 Q2
-6 -20 8 -12
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 21 0
1 U
6901 0 0
2
44326.5 59
0
6 74112~
219 1976 759 0 7 32
0 3 16 27 16 14 115 26
0
0 0 4704 0
5 74112
4 -60 39 -52
2 Q3
-6 -20 8 -12
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 21 0
1 U
842 0 0
2
44326.5 60
0
6 74112~
219 956 915 0 7 32
0 5 12 13 12 3 116 8
0
0 0 4704 0
5 74112
4 -60 39 -52
2 Q3
-7 -22 7 -14
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 23 0
1 U
3277 0 0
2
44326.5 61
0
8 4-In OR~
219 716 761 0 5 22
0 11 10 9 8 31
0
0 0 96 180
4 4072
-14 -24 14 -16
4 U18A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 24 0
1 U
4212 0 0
2
44326.5 62
0
9 2-In AND~
219 1639 772 0 3 22
0 6 7 14
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 20 0
1 U
4720 0 0
2
44326.5 63
0
9 2-In AND~
219 958 819 0 3 22
0 6 7 5
0
0 0 96 270
6 74LS08
-21 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 20 0
1 U
5551 0 0
2
44326.5 64
0
7 Pulser~
4 87 1104 0 10 12
0 117 118 15 4 0 0 5 5 5
7
0
0 0 4640 0
0
3 CLK
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6986 0 0
2
44326.5 65
0
260
3 0 2 0 0 4096 0 1 0 0 210 3
133 440
91 440
91 481
2 0 3 0 0 4096 3 1 0 0 114 2
133 426
115 426
0 4 4 0 0 8320 0 0 67 96 0 3
1020 958
1020 1104
117 1104
5 0 5 0 0 8192 0 57 0 0 9 3
802 932
802 933
883 933
3 1 5 0 0 0 0 66 63 0 0 2
956 842
956 852
1 0 3 0 0 12288 3 58 0 0 7 5
883 854
883 768
993 768
993 934
956 934
5 0 3 0 0 0 3 63 0 0 179 2
956 927
956 1056
0 1 3 0 0 0 3 0 56 13 0 3
803 854
803 855
717 855
0 5 5 0 0 8320 0 0 58 5 0 5
956 843
918 843
918 933
883 933
883 929
5 5 5 0 0 0 0 57 56 0 0 4
802 932
802 933
717 933
717 930
1 0 6 0 0 8192 0 66 0 0 206 5
965 797
965 787
661 787
661 608
611 608
0 2 7 0 0 8192 0 0 66 180 0 4
663 1065
663 794
947 794
947 797
1 1 3 0 0 0 3 58 57 0 0 3
883 854
802 854
802 857
4 7 8 0 0 4224 0 64 63 0 0 5
739 747
982 747
982 880
980 880
980 879
3 7 9 0 0 4224 0 64 58 0 0 5
739 756
912 756
912 880
907 880
907 881
2 7 10 0 0 8320 0 64 57 0 0 5
739 765
835 765
835 883
826 883
826 884
7 1 11 0 0 8320 0 56 64 0 0 4
741 882
752 882
752 774
739 774
0 4 12 0 0 4096 0 0 63 19 0 3
923 880
923 897
932 897
0 2 12 0 0 8192 0 0 63 46 0 6
846 800
923 800
923 880
935 880
935 879
932 879
6 3 13 0 0 8320 0 58 63 0 0 4
913 899
916 899
916 888
926 888
4 0 12 0 0 0 0 56 0 0 45 3
693 900
680 900
680 882
0 0 12 0 0 0 0 0 0 45 153 3
679 801
679 799
678 799
0 1 6 0 0 4224 0 0 65 62 0 4
593 414
1610 414
1610 763
1615 763
2 4 7 0 0 0 0 65 11 0 0 3
1615 781
1557 781
1557 772
5 3 14 0 0 4224 0 59 65 0 0 2
1749 772
1660 772
0 3 15 0 0 4224 0 0 59 29 0 4
670 1094
1688 1094
1688 733
1719 733
2 0 12 0 0 0 0 58 0 0 46 2
859 881
846 881
2 0 12 0 0 0 0 57 0 0 45 2
778 884
765 884
3 0 15 0 0 0 0 56 0 0 196 4
687 891
670 891
670 1095
511 1095
3 0 15 0 0 0 0 20 0 0 196 2
520 1021
513 1021
3 0 15 0 0 0 0 19 0 0 196 2
520 919
513 919
1 1 3 0 0 0 3 61 62 0 0 4
1899 696
1899 697
1976 697
1976 696
5 5 14 0 0 0 0 61 62 0 0 4
1899 771
1899 772
1976 772
1976 771
4 0 16 0 0 4096 0 62 0 0 63 2
1952 741
1942 741
4 0 16 0 0 0 0 61 0 0 64 2
1875 741
1866 741
5 5 14 0 0 0 0 61 60 0 0 4
1899 771
1899 772
1827 772
1827 771
5 5 14 0 0 0 0 60 59 0 0 3
1827 771
1827 772
1749 772
1 1 3 0 0 0 3 61 60 0 0 4
1899 696
1899 697
1827 697
1827 696
1 1 3 0 0 0 3 60 59 0 0 3
1827 696
1827 697
1749 697
4 0 16 0 0 0 0 60 0 0 65 5
1803 741
1803 740
1799 740
1799 741
1795 741
7 0 17 0 0 0 0 60 0 0 60 2
1851 723
1851 723
4 0 16 0 0 0 0 59 0 0 66 2
1725 742
1715 742
3 6 18 0 0 4224 0 58 57 0 0 4
853 890
840 890
840 902
832 902
3 6 19 0 0 4224 0 57 56 0 0 4
772 893
756 893
756 900
747 900
2 4 12 0 0 32768 0 56 57 0 0 10
693 882
679 882
679 883
680 883
680 823
679 823
679 800
765 800
765 902
778 902
0 4 12 0 0 0 0 0 58 45 0 4
764 800
846 800
846 899
859 899
12 11 20 0 0 4096 0 55 0 0 220 2
1918 558
1918 395
11 10 21 0 0 4096 0 55 0 0 220 2
1900 558
1900 395
10 9 22 0 0 4096 0 55 0 0 220 2
1882 558
1882 395
9 8 23 0 0 4096 0 55 0 0 220 2
1864 558
1864 395
3 3 15 0 0 0 0 20 20 0 0 2
520 1021
520 1021
3 0 4 0 0 0 0 2 0 0 116 5
1031 742
959 742
959 406
467 406
467 348
0 1 24 0 0 12288 0 0 34 202 0 4
603 444
801 444
801 155
511 155
5 1 25 0 0 12416 0 20 55 0 0 6
574 1021
603 1021
603 1073
1666 1073
1666 628
1855 628
5 7 25 0 0 0 0 55 55 0 0 2
1891 628
1909 628
3 5 25 0 0 0 0 55 55 0 0 2
1873 628
1891 628
1 3 25 0 0 0 0 55 55 0 0 2
1855 628
1873 628
8 7 26 0 0 8320 0 55 62 0 0 5
1918 622
1918 638
2011 638
2011 723
2000 723
6 0 27 0 0 12416 0 55 0 0 67 4
1900 622
1900 645
1928 645
1928 723
4 0 17 0 0 12416 0 55 0 0 68 4
1882 622
1882 646
1851 646
1851 723
2 0 28 0 0 12416 0 55 0 0 69 4
1864 622
1864 638
1787 638
1787 723
0 17 6 0 0 0 0 0 32 206 0 5
593 608
593 414
265 414
265 308
237 308
2 0 16 0 0 12288 0 62 0 0 64 4
1952 723
1942 723
1942 779
1865 779
0 2 16 0 0 0 0 0 61 65 0 4
1795 779
1866 779
1866 723
1875 723
2 0 16 0 0 12288 0 60 0 0 66 4
1803 723
1795 723
1795 779
1715 779
0 2 16 0 0 12416 0 0 59 75 0 6
581 901
621 901
621 1084
1715 1084
1715 724
1725 724
7 3 27 0 0 0 0 61 62 0 0 4
1923 723
1936 723
1936 732
1946 732
0 3 17 0 0 0 0 0 61 0 0 4
1845 723
1861 723
1861 732
1869 732
7 3 28 0 0 0 0 59 60 0 0 6
1773 724
1787 724
1787 723
1787 723
1787 732
1797 732
0 1 3 0 0 4096 3 0 11 39 0 2
1749 697
1557 697
0 1 29 0 0 8192 0 0 52 84 0 3
422 808
379 808
379 970
2 0 30 0 0 4096 0 52 0 0 73 2
379 988
351 988
2 1 30 0 0 8320 0 54 53 0 0 5
650 844
650 959
351 959
351 1018
381 1018
1 0 31 0 0 4096 0 54 0 0 86 2
650 808
650 761
0 2 16 0 0 0 0 0 53 87 0 5
581 901
581 955
345 955
345 1036
381 1036
2 3 32 0 0 8320 0 51 53 0 0 4
444 1012
435 1012
435 1027
426 1027
1 3 33 0 0 8320 0 51 52 0 0 4
444 994
435 994
435 979
424 979
2 3 34 0 0 4224 0 20 51 0 0 2
520 1003
490 1003
0 1 35 0 0 4096 0 0 50 89 0 3
345 754
345 911
389 911
2 2 36 0 0 8320 0 49 50 0 0 3
444 910
444 911
425 911
1 0 12 0 0 12288 0 49 0 0 90 5
444 892
433 892
433 855
596 855
596 798
2 3 37 0 0 4224 0 19 49 0 0 2
520 901
489 901
0 1 31 0 0 0 0 0 48 86 0 3
435 761
435 790
445 790
0 2 29 0 0 8192 0 0 48 101 0 5
597 696
597 748
422 748
422 808
445 808
2 3 38 0 0 4224 0 18 48 0 0 2
521 799
490 799
5 2 31 0 0 4224 0 64 47 0 0 4
689 761
371 761
371 743
376 743
6 1 16 0 0 0 0 19 47 0 0 6
568 901
581 901
581 863
362 863
362 725
376 725
3 3 39 0 0 8320 0 47 45 0 0 4
421 734
432 734
432 705
442 705
5 1 35 0 0 12416 0 42 46 0 0 8
1585 924
1593 924
1593 986
637 986
637 754
345 754
345 687
377 687
0 2 12 0 0 8192 0 0 46 153 0 5
596 799
596 766
354 766
354 705
377 705
3 2 40 0 0 4224 0 46 45 0 0 2
422 696
443 696
0 1 41 0 0 8192 0 0 45 157 0 5
617 590
617 648
432 648
432 687
442 687
2 4 42 0 0 4224 0 17 45 0 0 2
522 696
488 696
1 0 3 0 0 8192 3 42 0 0 179 3
1555 879
1555 848
1008 848
4 0 7 0 0 8192 0 42 0 0 180 3
1555 954
1555 967
1055 967
0 3 4 0 0 0 0 0 42 164 0 5
1020 778
1020 959
1514 959
1514 924
1531 924
2 6 43 0 0 8320 0 41 42 0 0 5
1393 946
1393 971
1601 971
1601 906
1579 906
6 1 44 0 0 12416 0 11 40 0 0 5
1581 724
1596 724
1596 843
1393 843
1393 865
2 1 45 0 0 4224 0 44 41 0 0 2
1329 928
1393 928
1 0 29 0 0 0 0 44 0 0 101 3
1293 928
1257 928
1257 883
6 2 29 0 0 4224 0 17 40 0 0 4
570 696
999 696
999 883
1393 883
2 3 46 0 0 8320 0 42 43 0 0 3
1531 906
1531 905
1512 905
3 2 47 0 0 8320 0 41 43 0 0 4
1438 937
1456 937
1456 914
1466 914
3 1 48 0 0 8320 0 40 43 0 0 4
1438 874
1456 874
1456 896
1466 896
6 4 49 0 0 12416 0 38 39 0 0 5
550 284
562 284
562 376
381 376
381 300
6 3 50 0 0 12416 0 37 39 0 0 5
623 283
633 283
633 372
387 372
387 300
6 2 51 0 0 12416 0 36 39 0 0 5
693 283
704 283
704 366
393 366
393 300
6 1 52 0 0 12416 0 35 39 0 0 5
766 283
789 283
789 361
399 361
399 300
2 8 23 0 0 12416 0 34 0 0 220 4
502 155
502 110
311 110
311 395
4 9 22 0 0 12416 0 34 0 0 220 4
484 155
484 115
323 115
323 395
6 10 21 0 0 12416 0 34 0 0 220 4
466 155
466 121
335 121
335 395
8 11 20 0 0 12416 0 34 0 0 220 4
448 155
448 127
346 127
346 395
0 0 7 0 0 0 0 0 0 120 192 2
526 337
526 426
0 1 3 0 0 0 3 0 38 186 0 6
92 583
115 583
115 404
462 404
462 257
526 257
0 3 4 0 0 0 0 0 37 117 0 4
637 348
566 348
566 301
575 301
3 0 4 0 0 0 0 38 0 0 115 4
502 302
467 302
467 348
566 348
3 3 4 0 0 0 0 36 35 0 0 6
645 301
637 301
637 348
708 348
708 301
718 301
0 4 7 0 0 0 0 0 35 119 0 3
668 337
742 337
742 331
0 4 7 0 0 0 0 0 36 120 0 3
599 337
669 337
669 331
4 4 7 0 0 0 0 38 37 0 0 4
526 332
526 337
599 337
599 331
1 1 3 0 0 0 3 36 35 0 0 4
669 256
669 257
742 257
742 256
1 1 3 0 0 0 3 37 36 0 0 4
599 256
599 257
669 257
669 256
1 1 3 0 0 0 3 38 37 0 0 3
526 257
599 257
599 256
6 3 52 0 0 0 0 35 34 0 0 4
766 283
766 136
493 136
493 155
6 5 51 0 0 0 0 36 34 0 0 4
693 283
693 141
475 141
475 155
6 7 50 0 0 0 0 37 34 0 0 4
623 283
623 145
457 145
457 155
6 9 49 0 0 0 0 38 34 0 0 4
550 284
550 149
439 149
439 155
1 10 2 0 0 0 0 33 34 0 0 4
430 149
430 146
430 146
430 149
11 2 53 0 0 8320 0 34 35 0 0 5
493 219
493 222
708 222
708 283
718 283
12 2 54 0 0 8320 0 34 36 0 0 5
475 219
475 227
637 227
637 283
645 283
13 2 55 0 0 8320 0 34 37 0 0 5
457 219
457 233
566 233
566 283
575 283
14 2 56 0 0 4224 0 34 38 0 0 3
439 219
439 284
502 284
17 18 6 0 0 0 0 32 32 0 0 2
237 308
192 308
9 0 57 0 0 4096 0 32 0 0 220 2
228 378
228 395
10 1 58 0 0 4096 0 32 0 0 220 2
219 378
219 395
11 2 59 0 0 4096 0 32 0 0 220 2
210 378
210 395
12 3 60 0 0 4096 0 32 0 0 220 2
201 378
201 395
13 4 61 0 0 4096 0 32 0 0 220 2
183 378
183 395
14 5 62 0 0 4096 0 32 0 0 220 2
174 378
174 395
15 6 63 0 0 4096 0 32 0 0 220 2
165 378
165 395
16 7 64 0 0 4096 0 32 0 0 220 2
156 378
156 395
1 1 65 0 0 8320 0 31 32 0 0 3
224 299
228 299
228 314
2 2 66 0 0 4224 0 32 31 0 0 3
219 314
219 299
218 299
3 3 67 0 0 4224 0 32 31 0 0 3
210 314
210 299
212 299
4 4 68 0 0 4224 0 32 31 0 0 3
201 314
201 299
206 299
1 5 69 0 0 8320 0 30 32 0 0 3
178 300
183 300
183 314
2 6 70 0 0 8320 0 30 32 0 0 3
172 300
174 300
174 314
3 7 71 0 0 8320 0 30 32 0 0 3
166 300
165 300
165 314
4 8 72 0 0 8320 0 30 32 0 0 3
160 300
156 300
156 314
0 12 12 0 0 0 0 0 9 151 0 3
1320 609
1460 609
1460 617
0 12 12 0 0 0 0 0 10 152 0 3
1174 609
1321 609
1321 617
0 12 12 0 0 0 0 0 8 153 0 3
1035 609
1175 609
1175 618
6 12 12 0 0 12416 0 18 7 0 0 5
569 799
678 799
678 609
1036 609
1036 618
11 0 41 0 0 0 0 9 0 0 155 3
1469 617
1469 590
1330 590
11 0 41 0 0 0 0 10 0 0 156 3
1330 617
1330 590
1184 590
11 0 41 0 0 0 0 8 0 0 157 3
1184 618
1184 590
1045 590
11 6 41 0 0 8320 0 7 16 0 0 3
1045 618
1045 590
572 590
3 0 4 0 0 0 0 11 0 0 159 4
1533 742
1521 742
1521 778
1452 778
3 0 4 0 0 0 0 12 0 0 160 4
1460 742
1452 742
1452 778
1383 778
3 0 4 0 0 0 0 13 0 0 161 4
1390 742
1383 742
1383 778
1305 778
3 0 4 0 0 0 0 14 0 0 162 4
1316 742
1305 742
1305 778
1236 778
3 0 4 0 0 0 0 5 0 0 163 4
1247 742
1236 742
1236 778
1167 778
3 0 4 0 0 0 0 4 0 0 164 4
1175 742
1167 742
1167 778
1105 778
3 0 4 0 0 0 0 3 0 0 52 4
1105 742
1105 778
1020 778
1020 742
4 4 7 0 0 0 0 12 11 0 0 2
1484 772
1557 772
4 4 7 0 0 0 0 12 13 0 0 2
1484 772
1414 772
4 4 7 0 0 0 0 14 13 0 0 2
1340 772
1414 772
4 4 7 0 0 0 0 5 14 0 0 2
1271 772
1340 772
4 4 7 0 0 0 0 4 5 0 0 2
1199 772
1271 772
4 4 7 0 0 0 0 3 4 0 0 2
1129 772
1199 772
4 4 7 0 0 0 0 3 2 0 0 2
1129 772
1055 772
1 1 3 0 0 0 3 12 11 0 0 2
1484 697
1557 697
1 1 3 0 0 0 3 13 12 0 0 2
1414 697
1484 697
1 1 3 0 0 0 3 14 13 0 0 2
1340 697
1414 697
1 1 3 0 0 0 3 5 14 0 0 2
1271 697
1340 697
1 1 3 0 0 0 3 4 5 0 0 2
1199 697
1271 697
1 1 3 0 0 0 3 3 4 0 0 2
1129 697
1199 697
1 1 3 0 0 0 3 2 3 0 0 2
1055 697
1129 697
0 1 3 0 0 8320 3 0 2 186 0 5
92 669
92 1056
1008 1056
1008 697
1055 697
0 4 7 0 0 8320 0 0 2 207 0 4
184 560
184 1065
1055 1065
1055 772
1 0 3 0 0 0 3 20 0 0 182 3
544 976
587 976
587 874
1 0 3 0 0 0 3 19 0 0 183 3
544 874
587 874
587 772
1 0 3 0 0 0 3 18 0 0 185 3
545 772
587 772
587 669
1 4 3 0 0 0 3 16 15 0 0 2
548 563
548 538
1 1 3 0 0 0 3 17 16 0 0 5
546 669
587 669
587 558
548 558
548 563
1 1 3 0 0 0 3 29 17 0 0 3
92 564
92 669
546 669
0 4 7 0 0 0 0 0 20 188 0 3
505 948
505 1051
544 1051
0 4 7 0 0 0 0 0 19 189 0 3
505 846
505 949
544 949
0 4 7 0 0 0 0 0 18 190 0 3
505 743
505 847
545 847
0 4 7 0 0 0 0 0 17 191 0 3
505 638
505 744
546 744
4 0 7 0 0 0 0 16 0 0 192 4
548 638
505 638
505 451
548 451
1 0 7 0 0 0 0 15 0 0 207 3
548 463
548 426
183 426
0 3 15 0 0 0 0 0 15 194 0 3
513 609
513 508
524 508
0 3 15 0 0 0 0 0 16 195 0 3
513 714
513 608
524 608
0 3 15 0 0 0 0 0 17 196 0 3
513 817
513 714
522 714
3 3 15 0 0 0 0 67 18 0 0 4
111 1095
513 1095
513 817
521 817
2 3 73 0 0 4224 0 16 27 0 0 2
524 590
492 590
1 0 74 0 0 8192 0 27 0 0 204 3
447 581
432 581
432 550
0 2 75 0 0 12288 0 0 27 208 0 4
325 522
365 522
365 599
447 599
2 1 76 0 0 4224 0 28 26 0 0 2
369 490
375 490
1 0 75 0 0 0 0 28 0 0 208 2
333 490
325 490
6 1 24 0 0 8320 0 20 25 0 0 6
568 1003
603 1003
603 444
439 444
439 481
447 481
3 2 77 0 0 4224 0 25 15 0 0 2
493 490
524 490
6 2 74 0 0 12416 0 15 26 0 0 5
572 490
612 490
612 550
375 550
375 508
2 3 78 0 0 4224 0 25 26 0 0 2
447 499
420 499
5 3 6 0 0 0 0 16 24 0 0 6
578 608
612 608
612 656
229 656
229 569
243 569
1 2 7 0 0 0 0 1 24 0 0 4
172 426
184 426
184 560
243 560
3 1 75 0 0 12416 0 22 24 0 0 6
293 490
325 490
325 522
229 522
229 551
243 551
4 2 79 0 0 12416 0 24 22 0 0 6
294 560
325 560
325 530
235 530
235 499
242 499
2 1 2 0 0 4096 0 21 23 0 0 3
135 481
91 481
91 512
1 1 80 0 0 4224 0 21 22 0 0 2
169 481
242 481
2 0 57 0 0 4224 0 9 0 0 220 2
1550 617
1550 395
7 1 58 0 0 4224 0 9 0 0 220 2
1505 617
1505 395
2 2 59 0 0 4224 0 10 0 0 220 2
1411 617
1411 395
7 3 60 0 0 4224 0 10 0 0 220 2
1366 617
1366 395
2 4 61 0 0 4224 0 8 0 0 220 2
1265 618
1265 395
7 5 62 0 0 4224 0 8 0 0 220 2
1220 618
1220 395
2 6 63 0 0 4224 0 7 0 0 220 2
1126 618
1126 395
7 7 64 0 0 4224 0 7 0 0 220 2
1081 618
1081 395
-215140 0 1 0 0 4256 0 0 0 0 0 2
75 395
2065 395
3 0 81 0 0 8192 0 9 0 0 231 3
1541 617
1541 602
1514 602
8 0 82 0 0 8192 0 9 0 0 234 3
1496 617
1496 602
1442 602
3 0 83 0 0 8192 0 10 0 0 235 3
1402 617
1402 602
1375 602
8 0 84 0 0 8192 0 10 0 0 246 3
1357 617
1357 602
1295 602
3 0 85 0 0 8192 0 8 0 0 247 3
1256 618
1256 602
1229 602
8 0 86 0 0 8192 0 8 0 0 250 3
1211 618
1211 602
1157 602
8 0 2 0 0 0 0 7 0 0 255 2
1072 618
1072 575
3 0 87 0 0 8192 0 7 0 0 251 3
1117 618
1117 602
1090 602
1 0 44 0 0 0 0 9 0 0 230 2
1559 617
1559 583
6 4 44 0 0 0 0 11 9 0 0 4
1581 724
1581 583
1532 583
1532 617
0 6 81 0 0 8192 0 0 9 232 0 3
1485 583
1514 583
1514 617
6 9 81 0 0 12416 0 12 9 0 0 6
1508 724
1508 688
1447 688
1447 583
1487 583
1487 617
1 0 82 0 0 0 0 10 0 0 234 2
1420 617
1420 583
6 4 82 0 0 8320 0 13 10 0 0 5
1438 724
1442 724
1442 583
1393 583
1393 617
0 6 83 0 0 8192 0 0 10 236 0 3
1348 583
1375 583
1375 617
6 9 83 0 0 12416 0 14 10 0 0 6
1364 724
1364 688
1308 688
1308 583
1348 583
1348 617
5 0 2 0 0 8192 0 9 0 0 238 3
1523 611
1523 574
1478 574
10 0 2 0 0 8192 0 9 0 0 239 3
1478 611
1478 574
1384 574
5 0 2 0 0 0 0 10 0 0 240 4
1384 611
1384 574
1339 574
1339 575
10 0 2 0 0 8320 0 10 0 0 253 3
1339 611
1339 575
1238 575
14 2 88 0 0 12416 0 9 11 0 0 5
1541 681
1541 684
1521 684
1521 724
1533 724
13 2 89 0 0 8320 0 9 12 0 0 5
1496 681
1496 684
1452 684
1452 724
1460 724
14 2 90 0 0 12416 0 10 13 0 0 5
1402 681
1402 686
1383 686
1383 724
1390 724
13 2 91 0 0 8320 0 10 14 0 0 5
1357 681
1357 684
1305 684
1305 724
1316 724
1 0 84 0 0 0 0 8 0 0 246 2
1274 618
1274 584
6 4 84 0 0 4224 0 5 8 0 0 4
1295 724
1295 584
1247 584
1247 618
0 6 85 0 0 8192 0 0 8 248 0 3
1200 584
1229 584
1229 618
6 9 85 0 0 12416 0 4 8 0 0 6
1223 724
1223 689
1162 689
1162 584
1202 584
1202 618
1 0 86 0 0 0 0 7 0 0 250 2
1135 618
1135 584
6 4 86 0 0 8320 0 3 7 0 0 5
1153 724
1157 724
1157 584
1108 584
1108 618
0 6 87 0 0 8192 0 0 7 252 0 3
1063 584
1090 584
1090 618
6 9 87 0 0 12416 0 2 7 0 0 6
1079 724
1079 689
1023 689
1023 584
1063 584
1063 618
5 0 2 0 0 0 0 8 0 0 254 3
1238 612
1238 575
1193 575
10 0 2 0 0 0 0 8 0 0 255 3
1193 612
1193 575
1099 575
5 0 2 0 0 0 0 7 0 0 256 3
1099 612
1099 575
1054 575
10 1 2 0 0 0 0 7 6 0 0 3
1054 612
1054 575
973 575
14 2 92 0 0 12416 0 8 5 0 0 5
1256 682
1256 685
1236 685
1236 724
1247 724
13 2 93 0 0 8320 0 8 4 0 0 5
1211 682
1211 685
1167 685
1167 724
1175 724
14 2 94 0 0 12416 0 7 3 0 0 5
1117 682
1117 687
1098 687
1098 724
1105 724
13 2 95 0 0 8320 0 7 2 0 0 5
1072 682
1072 685
1020 685
1020 724
1031 724
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
1830 778 2002 797
1847 792 1984 805
17 RIPPLE UP COUNTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
701 935 936 954
718 949 918 962
25 MOD-8 RIPPLE DOWN COUNTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 44
898 9 1261 33
903 13 1255 29
44 NUMBER OF ONES IN BINARY BIT PATTERN COUNTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
146 207 237 231
151 211 231 227
10 INPUT UNIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
860 608 911 632
865 612 905 628
5 SHIFT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1269 540 1360 564
1274 544 1354 560
10 REGISTER R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
861 567 904 591
866 571 898 587
4 LOAD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
546 162 701 186
551 166 695 182
18 1's COUNT REGISTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
354 221 437 245
359 225 431 241
9 1's COUNT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
453 73 552 97
458 77 546 93
11 OUTPUT UNIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
343 1057 475 1076
360 1071 457 1084
12 CONTROL UNIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
1260 448 1367 467
1277 462 1349 475
9 DATA UNIT
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
